library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity plane_rom is
	Port (address : in STD_LOGIC_VECTOR(9 downto 0);
		   data_out : out STD_LOGIC_VECTOR(11 downto 0));
end plane_rom;

architecture Behavioral of plane_rom is
	type ROM_Type is array (0 to 199) of STD_LOGIC_VECTOR(11 downto 0);
	constant ROM : ROM_Type := (
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"010001000101",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"010001000101",
		"010001000101",
		"010001000101",
		"011001000011",
		"011001000011",
		"000000000000",
		"011001000011",
		"010001000101",
		"010001000101",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"011001000011",
		"011001000011",
		"010001000101",
		"010001000101",
		"011001000011",
		"000000000000",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"011001000011",
		"010001000101",
		"011001000011",
		"011001000011",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"011001000011",
		"000000000000",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"011001000011",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"011001000011",
		"111111101100",
		"111111101100",
		"111111101100",
		"010001000101",
		"010001000101",
		"010001000101",
		"011001000011",
		"011001000011",
		"111111101100",
		"111111101100",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"010001000101",
		"010001000101",
		"010001000101",
		"010001000101",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"011001000011",
		"011001000011",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"011001000011",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"011001000011",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"111111101100",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"011001000011",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000",
		"000000000000"
	);
begin
	process(address)
	begin
		data_out <= ROM(to_integer(unsigned(address)));
	end process;
end Behavioral;
